-- converted by jbboot_bin2vhdl.py
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity jbboot is
   port
   (
        clk: in std_logic;
        addr: in std_logic_vector(9 downto 0);
        data: out std_logic_vector(15 downto 0)
   );
end jbboot;

architecture arch of jbboot is
   type rom_type is array (0 to 1023) of std_logic_vector(15 downto 0);
   constant rom_data: rom_type := (
x"0001",x"0000",x"0000",x"0008",x"4df9",x"00df",x"f000",x"3d7c",
x"9000",x"0100",x"3d7c",x"0000",x"0102",x"3d7c",x"0000",x"0104",
x"3d7c",x"0000",x"0108",x"3d7c",x"0000",x"010a",x"6100",x"02de",
x"3d7c",x"003c",x"0092",x"3d7c",x"00d4",x"0094",x"3d7c",x"2c81",
x"008e",x"3d7c",x"f4c1",x"0090",x"3d7c",x"037f",x"0180",x"3d7c",
x"0fff",x"0182",x"41fa",x"02d2",x"43f9",x"0000",x"c100",x"7002",
x"22d8",x"4e71",x"51c8",x"fffa",x"2d7c",x"0000",x"c100",x"0080",
x"3d40",x"0088",x"3d7c",x"8390",x"0096",x"3d7c",x"7fff",x"009e",
x"41fa",x"064b",x"6100",x"025e",x"41fa",x"06e3",x"6100",x"0256",
x"41fa",x"06f5",x"6100",x"024e",x"41fa",x"059a",x"6100",x"0246",
x"302e",x"0004",x"e048",x"0200",x"007f",x"6100",x"01d0",x"41fa",
x"0592",x"0801",x"0004",x"6704",x"41fa",x"058f",x"6100",x"0226",
x"41fa",x"058f",x"6100",x"021e",x"302e",x"007c",x"6100",x"01ae",
x"700a",x"6100",x"01c0",x"700a",x"6100",x"01ba",x"13fc",x"0003",
x"00bf",x"e201",x"13fc",x"0000",x"00bf",x"e001",x"13fc",x"00ff",
x"00bf",x"d300",x"13fc",x"00f7",x"00bf",x"d100",x"13fc",x"00f6",
x"00bf",x"d100",x"13fc",x"00f7",x"00bf",x"d100",x"0839",x"0002",
x"00bf",x"e001",x"67e6",x"303c",x"000c",x"6100",x"0128",x"307c",
x"4000",x"0c58",x"aaca",x"6600",x"0108",x"3018",x"b07c",x"0001",
x"6626",x"2018",x"6100",x"010e",x"41f8",x"4000",x"0c10",x"00fe",
x"6608",x"3d7c",x"0f00",x"0180",x"5248",x"6100",x"0198",x"700a",
x"6100",x"0142",x"6000",x"00ea",x"b07c",x"0002",x"6600",x"0092",
x"2858",x"2a4c",x"2818",x"2a04",x"41fa",x"04f5",x"6100",x"0176",
x"200c",x"6100",x"00f8",x"41fa",x"04f6",x"6100",x"0168",x"2004",
x"6100",x"00ea",x"700a",x"6100",x"010c",x"41fa",x"04ec",x"6100",
x"0154",x"947c",x"0021",x"47eb",x"ffdf",x"2c05",x"ea8e",x"bc84",
x"6d02",x"2c04",x"3006",x"6100",x"009c",x"3006",x"e448",x"5340",
x"28d8",x"4e71",x"51c8",x"fffa",x"707f",x"6100",x"00d8",x"0879",
x"0001",x"00bf",x"e001",x"9886",x"6ed0",x"bbfc",x"00f8",x"0000",
x"6616",x"babc",x"0004",x"0000",x"660e",x"284d",x"d9c5",x"7aff",
x"28dd",x"4e71",x"51cd",x"fffa",x"700a",x"6100",x"00a8",x"6050",
x"b07c",x"0003",x"6610",x"08f9",x"0001",x"00bf",x"e001",x"4a39",
x"00bf",x"c000",x"60fe",x"b07c",x"0004",x"660e",x"2858",x"2818",
x"7000",x"28c0",x"5984",x"6efa",x"6026",x"3e00",x"3d7c",x"0f00",
x"0180",x"41fa",x"0495",x"6100",x"00bc",x"3007",x"6146",x"60fe",
x"3d7c",x"0f00",x"0180",x"41fa",x"0463",x"6100",x"00a8",x"60ee",
x"6000",x"fed4",x"3d7c",x"0002",x"009c",x"307c",x"4000",x"2d48",
x"0020",x"e248",x"0040",x"8000",x"3d40",x"0024",x"3d40",x"0024",
x"302e",x"001e",x"0800",x"0001",x"67f6",x"4e75",x"4840",x"6104",
x"4841",x"2001",x"e058",x"6104",x"2001",x"e058",x"2200",x"e808",
x"6106",x"2001",x"0200",x"000f",x"d03c",x"0030",x"b03c",x"0039",
x"6f02",x"5e00",x"224b",x"528b",x"b03c",x"000a",x"660c",x"96c2",
x"343c",x"0000",x"47eb",x"027f",x"6028",x"4880",x"907c",x"0020",
x"e740",x"41fa",x"0080",x"d0c0",x"7007",x"1298",x"43e9",x"0050",
x"51c8",x"fff8",x"5242",x"b47c",x"0050",x"6616",x"7400",x"47eb",
x"0230",x"5243",x"b67c",x"0019",x"6608",x"5343",x"47eb",x"fd80",
x"6112",x"4e75",x"2448",x"224b",x"7000",x"101a",x"6704",x"61a4",
x"60f4",x"4e75",x"41f9",x"0000",x"8000",x"43e8",x"0280",x"303c",
x"0f9f",x"20d9",x"4e71",x"51c8",x"fffa",x"4e75",x"7400",x"7600",
x"47f9",x"0000",x"8000",x"204b",x"7000",x"323c",x"103f",x"20c0",
x"4e71",x"51c9",x"fffa",x"4e75",x"00e0",x"0000",x"00e2",x"8000",
x"ffff",x"fffe",x"0000",x"0000",x"0000",x"0000",x"1818",x"1818",
x"1800",x"1800",x"6c6c",x"0000",x"0000",x"0000",x"6c6c",x"fe6c",
x"fe6c",x"6c00",x"183e",x"603c",x"067c",x"1800",x"0066",x"acd8",
x"366a",x"cc00",x"386c",x"6876",x"dcce",x"7b00",x"1818",x"3000",
x"0000",x"0000",x"0c18",x"3030",x"3018",x"0c00",x"3018",x"0c0c",
x"0c18",x"3000",x"0066",x"3cff",x"3c66",x"0000",x"0018",x"187e",
x"1818",x"0000",x"0000",x"0000",x"0018",x"1830",x"0000",x"007e",
x"0000",x"0000",x"0000",x"0000",x"0018",x"1800",x"0306",x"0c18",
x"3060",x"c000",x"3c66",x"6e7e",x"7666",x"3c00",x"1838",x"7818",
x"1818",x"1800",x"3c66",x"060c",x"1830",x"7e00",x"3c66",x"061c",
x"0666",x"3c00",x"1c3c",x"6ccc",x"fe0c",x"0c00",x"7e60",x"7c06",
x"0666",x"3c00",x"1c30",x"607c",x"6666",x"3c00",x"7e06",x"060c",
x"1818",x"1800",x"3c66",x"663c",x"6666",x"3c00",x"3c66",x"663e",
x"060c",x"3800",x"0018",x"1800",x"0018",x"1800",x"0018",x"1800",
x"0018",x"1830",x"0006",x"1860",x"1806",x"0000",x"0000",x"7e00",
x"7e00",x"0000",x"0060",x"1806",x"1860",x"0000",x"3c66",x"060c",
x"1800",x"1800",x"7cc6",x"ded6",x"dec0",x"7800",x"3c66",x"667e",
x"6666",x"6600",x"7c66",x"667c",x"6666",x"7c00",x"1e30",x"6060",
x"6030",x"1e00",x"786c",x"6666",x"666c",x"7800",x"7e60",x"6078",
x"6060",x"7e00",x"7e60",x"6078",x"6060",x"6000",x"3c66",x"606e",
x"6666",x"3e00",x"6666",x"667e",x"6666",x"6600",x"3c18",x"1818",
x"1818",x"3c00",x"0606",x"0606",x"0666",x"3c00",x"c6cc",x"d8f0",
x"d8cc",x"c600",x"6060",x"6060",x"6060",x"7e00",x"c6ee",x"fed6",
x"c6c6",x"c600",x"c6e6",x"f6de",x"cec6",x"c600",x"3c66",x"6666",
x"6666",x"3c00",x"7c66",x"667c",x"6060",x"6000",x"78cc",x"cccc",
x"ccdc",x"7e00",x"7c66",x"667c",x"6c66",x"6600",x"3c66",x"703c",
x"0e66",x"3c00",x"7e18",x"1818",x"1818",x"1800",x"6666",x"6666",
x"6666",x"3c00",x"6666",x"6666",x"3c3c",x"1800",x"c6c6",x"c6d6",
x"feee",x"c600",x"c366",x"3c18",x"3c66",x"c300",x"c366",x"3c18",
x"1818",x"1800",x"fe0c",x"1830",x"60c0",x"fe00",x"3c30",x"3030",
x"3030",x"3c00",x"c060",x"3018",x"0c06",x"0300",x"3c0c",x"0c0c",
x"0c0c",x"3c00",x"1038",x"6cc6",x"0000",x"0000",x"0000",x"0000",
x"0000",x"00fe",x"1818",x"0c00",x"0000",x"0000",x"0000",x"3c06",
x"3e66",x"3e00",x"6060",x"7c66",x"6666",x"7c00",x"0000",x"3c60",
x"6060",x"3c00",x"0606",x"3e66",x"6666",x"3e00",x"0000",x"3c66",
x"7e60",x"3c00",x"1c30",x"7c30",x"3030",x"3000",x"0000",x"3e66",
x"663e",x"063c",x"6060",x"7c66",x"6666",x"6600",x"1800",x"1818",
x"1818",x"0c00",x"0c00",x"0c0c",x"0c0c",x"0c78",x"6060",x"666c",
x"786c",x"6600",x"1818",x"1818",x"1818",x"0c00",x"0000",x"ecfe",
x"d6c6",x"c600",x"0000",x"7c66",x"6666",x"6600",x"0000",x"3c66",
x"6666",x"3c00",x"0000",x"7c66",x"667c",x"6060",x"0000",x"3e66",
x"663e",x"0606",x"0000",x"7c66",x"6060",x"6000",x"0000",x"3c60",
x"3c06",x"7c00",x"3030",x"7c30",x"3030",x"1c00",x"0000",x"6666",
x"6666",x"3e00",x"0000",x"6666",x"663c",x"1800",x"0000",x"c6c6",
x"d6fe",x"6c00",x"0000",x"c66c",x"386c",x"c600",x"0000",x"6666",
x"663c",x"1830",x"0000",x"7e0c",x"1830",x"7e00",x"0e18",x"1870",
x"1818",x"0e00",x"1818",x"1818",x"1818",x"1800",x"7018",x"180e",
x"1818",x"7000",x"729c",x"0000",x"0000",x"0000",x"fefe",x"fefe",
x"fefe",x"fe00",x"0a0a",x"4167",x"6e75",x"7320",x"4944",x"3a20",
x"2400",x"2028",x"5041",x"4c29",x"0020",x"284e",x"5453",x"4329",
x"0020",x"4465",x"6e69",x"7365",x"2049",x"443a",x"2024",x"004d",
x"656d",x"6f72",x"7920",x"6261",x"7365",x"3a20",x"2400",x"2c20",
x"7369",x"7a65",x"3a20",x"2400",x"5b5f",x"5f5f",x"5f5f",x"5f5f",
x"5f5f",x"5f5f",x"5f5f",x"5f5f",x"5f5f",x"5f5f",x"5f5f",x"5f5f",
x"5f5f",x"5f5f",x"5f5f",x"5f5f",x"5f5d",x"000a",x"496e",x"636f",
x"6d70",x"6174",x"6962",x"6c65",x"204d",x"656e",x"7565",x"2066",
x"6972",x"6d77",x"6172",x"6521",x"000a",x"556e",x"6b6e",x"6f77",
x"6e20",x"636f",x"6d6d",x"616e",x"643a",x"2024",x"004d",x"696e",
x"696d",x"6967",x"2062",x"7920",x"4465",x"6e6e",x"6973",x"2076",
x"616e",x"2057",x"6565",x"7265",x"6e20",x"0a42",x"7567",x"2066",
x"6978",x"6573",x"2c20",x"6d6f",x"6473",x"2061",x"6e64",x"2065",
x"7874",x"656e",x"7369",x"6f6e",x"7320",x"6279",x"204a",x"616b",
x"7562",x"2042",x"6564",x"6e61",x"7273",x"6b69",x"2061",x"6e64",
x"2053",x"6173",x"6368",x"6120",x"426f",x"696e",x"6720",x"0a54",
x"4736",x"384b",x"2e43",x"2028",x"3638",x"3030",x"3020",x"4950",
x"2043",x"6f72",x"6529",x"2061",x"6e64",x"2043",x"6861",x"6d65",
x"6c65",x"6f6e",x"2050",x"6f72",x"7420",x"6279",x"2054",x"6f62",
x"6961",x"7320",x"4775",x"6265",x"6e65",x"720a",x"000a",x"426f",
x"6f74",x"6c6f",x"6164",x"6572",x"2020",x"2020",x"3230",x"3130",
x"2d30",x"392d",x"3130",x"000a",x"4d69",x"6e69",x"6d69",x"6720",
x"636f",x"7265",x"2020",x"3230",x"3131",x"2d30",x"342d",x"3130",
others => (others => '0'));
   signal R_data: std_logic_vector(15 downto 0);
   signal R_addr: std_logic_vector(9 downto 0);
begin
   process(clk)
   begin
      if rising_edge(clk) then
         R_data <= rom_data(to_integer(unsigned(addr)));
      end if;
   end process;
   data <= R_data;
end arch;
